module sign_extend(
output reg [31:0] sign_ext_imm,
input [15:0] imm);







endmodule
