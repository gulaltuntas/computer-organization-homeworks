module my_xor (output [31:0] y, input [31:0] a, input [31:0] b);
	
	xor xor1 (y[0], a[0], b[0]);
	xor xor2 (y[1], a[1], b[1]);
	xor xor3 (y[2], a[2], b[2]);
	xor xor4 (y[3], a[3], b[3]);
	xor xor5 (y[4], a[4], b[4]);
	xor xor6 (y[5], a[5], b[5]);
	xor xor7 (y[6], a[6], b[6]);
	xor xor8 (y[7], a[7], b[7]);
	xor xor9 (y[8], a[8], b[8]);
	xor xor10 (y[9], a[9], b[9]);
	xor xor11 (y[10], a[10], b[10]);
	xor xor12 (y[11], a[11], b[11]);
	xor xor13 (y[12], a[12], b[12]);
	xor xor14 (y[13], a[13], b[13]);
	xor xor15 (y[14], a[14], b[14]);
	xor xor16 (y[15], a[15], b[15]);
	xor xor17 (y[16], a[16], b[16]);
	xor xor18 (y[17], a[17], b[17]);
	xor xor19 (y[18], a[18], b[18]);
	xor xor20 (y[19], a[19], b[19]);
	xor xor21 (y[20], a[20], b[20]);
	xor xor22 (y[21], a[21], b[21]);
	xor xor23 (y[22], a[22], b[22]);
	xor xor24 (y[23], a[23], b[23]);
	xor xor25 (y[24], a[24], b[24]);
	xor xor26 (y[25], a[25], b[25]);
	xor xor27 (y[26], a[26], b[26]);
	xor xor28 (y[27], a[27], b[27]);
	xor xor29 (y[28], a[28], b[28]);
	xor xor30 (y[29], a[29], b[29]);
	xor xor31 (y[30], a[30], b[30]);
	xor xor32 (y[31], a[31], b[31]);

	



endmodule
