module my_nor (output [31:0] y, input [31:0] a, input [31:0] b);

	nor nor1 (y[0], a[0], b[0]);
	nor nor2 (y[1], a[1], b[1]);
	nor nor3 (y[2], a[2], b[2]);
	nor nor4 (y[3], a[3], b[3]);
	nor nor5 (y[4], a[4], b[4]);
	nor nor6 (y[5], a[5], b[5]);
	nor nor7 (y[6], a[6], b[6]);
	nor nor8 (y[7], a[7], b[7]);
	nor nor9 (y[8], a[8], b[8]);
	nor nor10 (y[9], a[9], b[9]);
	nor nor11 (y[10], a[10], b[10]);
	nor nor12 (y[11], a[11], b[11]);
	nor nor13 (y[12], a[12], b[12]);
	nor nor14 (y[13], a[13], b[13]);
	nor nor15 (y[14], a[14], b[14]);
	nor nor16 (y[15], a[15], b[15]);
	nor nor17 (y[16], a[16], b[16]);
	nor nor18 (y[17], a[17], b[17]);
	nor nor19 (y[18], a[18], b[18]);
	nor nor20 (y[19], a[19], b[19]);
	nor nor21 (y[20], a[20], b[20]);
	nor nor22 (y[21], a[21], b[21]);
	nor nor23 (y[22], a[22], b[22]);
	nor nor24 (y[23], a[23], b[23]);
	nor nor25 (y[24], a[24], b[24]);
	nor nor26 (y[25], a[25], b[25]);
	nor nor27 (y[26], a[26], b[26]);
	nor nor28 (y[27], a[27], b[27]);
	nor nor29 (y[28], a[28], b[28]);
	nor nor30 (y[29], a[29], b[29]);
	nor nor31 (y[30], a[30], b[30]);
	nor nor32 (y[31], a[31], b[31]);

endmodule
